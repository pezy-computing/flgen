module baz;
endmodule
