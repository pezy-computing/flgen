module bar;
endmodule
