module foo_lib;
endmodule
